library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity audio_gen is 
port (
    master_clock: in std_logic;
    clock_12_out: out std_logic:='0';
    ledr: OUT std_logic;
    keys: in std_logic_vector(3 downto 0); 
    aud_bk: out std_logic:='0';
    aud_dalr: out std_logic:='0';
    aud_data_out: out std_logic
);
end audio_gen; 

architecture gen of audio_gen is 
    signal clk_en: std_logic:='0';
    signal send_flag: std_logic:='0';
    signal index: integer range 0 to 23:=0;
    signal sample_index: integer range 0 to 999:=0;
    signal aud_idx: std_logic := '0';
    signal aud_out: std_logic_vector(23 downto 0):=(others=>'0');
    type BinArrray is array(0 to 999) of std_logic_vector(23 downto 0);
    
    -- 1046 C6
    -- 1000
    signal aud_out_sample: BinArrray :=("000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110101000"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010011000"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010011000"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110101000"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110101000"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000011111"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000011111"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110100111"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010011000"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011"
    ,"000000000010111100100010"
    ,"000000000011001010000000"
    ,"000000000011011001011000"
    ,"000000000011101010010111"
    ,"000000000011111100101101"
    ,"000000000100010000000011"
    ,"000000000100100100000110"
    ,"000000000100111000011111"
    ,"000000000101001100111001"
    ,"000000000101100000111100"
    ,"000000000101110100010010"
    ,"000000000110000110100111"
    ,"000000000110010111100111"
    ,"000000000110100110111111"
    ,"000000000110110100011101"
    ,"000000000110111111110100"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000111010011011010"
    ,"000000000111010100110000"
    ,"000000000111010011011010"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110111111110100"
    ,"000000000110110100011101"
    ,"000000000110100110111111"
    ,"000000000110010111100111"
    ,"000000000110000110101000"
    ,"000000000101110100010010"
    ,"000000000101100000111100"
    ,"000000000101001100111001"
    ,"000000000100111000100000"
    ,"000000000100100100000110"
    ,"000000000100010000000011"
    ,"000000000011111100101101"
    ,"000000000011101010010111"
    ,"000000000011011001011000"
    ,"000000000011001010000000"
    ,"000000000010111100100010"
    ,"000000000010110001001011"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000010011101100101"
    ,"000000000010011100010000"
    ,"000000000010011101100101"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000010110001001011");
    
    
    -- 1318 E6
    -- 5000 
    signal aud_out_sample1: BinArrray:=("000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110100111"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110100111"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110100111"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110101000"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110100111"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110100111"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010010111"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010010111"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000011111"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000100000"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100"
    ,"000000000111010011011010"
    ,"000000000110100110111111"
    ,"000000000101001100111001"
    ,"000000000011101010011000"
    ,"000000000010101000001001"
    ,"000000000010100001100100"
    ,"000000000011011001011000"
    ,"000000000100111000100000"
    ,"000000000110010111100111"
    ,"000000000111001111011011"
    ,"000000000111001000110110"
    ,"000000000110000110101000"
    ,"000000000100100100000110"
    ,"000000000011001010000000"
    ,"000000000010011101100101"
    ,"000000000010110001001011"
    ,"000000000011111100101101"
    ,"000000000101100000111100"
    ,"000000000110110100011101"
    ,"000000000111010100110000"
    ,"000000000110110100011101"
    ,"000000000101100000111100"
    ,"000000000011111100101101"
    ,"000000000010110001001011"
    ,"000000000010011101100101"
    ,"000000000011001010000000"
    ,"000000000100100100000110"
    ,"000000000110000110100111"
    ,"000000000111001000110110"
    ,"000000000111001111011011"
    ,"000000000110010111100111"
    ,"000000000100111000011111"
    ,"000000000011011001011000"
    ,"000000000010100001100100"
    ,"000000000010101000001001"
    ,"000000000011101010011000"
    ,"000000000101001100111001"
    ,"000000000110100110111111"
    ,"000000000111010011011010"
    ,"000000000110111111110100"
    ,"000000000101110100010010"
    ,"000000000100010000000011"
    ,"000000000010111100100010"
    ,"000000000010011100010000"
    ,"000000000010111100100010"
    ,"000000000100010000000011"
    ,"000000000101110100010010"
    ,"000000000110111111110100");

    -- 1568 G6
    -- 10000
    signal aud_out_sample2: BinArrray :=("000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110100111"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000011111"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000011111"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010010111"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110101000"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010011000"
    ,"000000000110100110111111"
    ,"000000000110111111110100"
    ,"000000000100010000000011"
    ,"000000000010011100010000"
    ,"000000000100010000000011"
    ,"000000000110111111110100"
    ,"000000000110100110111111"
    ,"000000000011101010011000"
    ,"000000000010100001100100"
    ,"000000000100111000100000"
    ,"000000000111001111011011"
    ,"000000000110000110101000"
    ,"000000000011001010000000"
    ,"000000000010110001001011"
    ,"000000000101100000111100"
    ,"000000000111010100110000"
    ,"000000000101100000111100"
    ,"000000000010110001001011"
    ,"000000000011001010000000"
    ,"000000000110000110100111"
    ,"000000000111001111011011"
    ,"000000000100111000100000"
    ,"000000000010100001100100"
    ,"000000000011101010010111"
    ,"000000000110100110111111"
    ,"000000000110111111110100");
    
    



    -- 1979.5 B6
    -- 15000
    signal aud_out_sample3: BinArrray:=("000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000011111"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000011111"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000"
    ,"000000000010101000001001"
    ,"000000000110100110111111"
    ,"000000000101110100010010"
    ,"000000000010011100010000"
    ,"000000000101110100010010"
    ,"000000000110100110111111"
    ,"000000000010101000001001"
    ,"000000000100111000100000"
    ,"000000000111001000110110"
    ,"000000000011001010000000"
    ,"000000000011111100101101"
    ,"000000000111010100110000"
    ,"000000000011111100101101"
    ,"000000000011001010000000"
    ,"000000000111001000110110"
    ,"000000000100111000100000");

    signal daclrc_count: integer range 0 to 519:=0;
    signal data_clock: std_logic:='0';
    signal aud_out_bit: std_logic;  
    constant ARRAY_SIZE: natural :=1000;
    signal bk_count: integer range 0 to 15:=0;
    signal aud_bk_clock: std_logic:='0';
    signal clock_12_count: integer range 0 to 1:=0;
    signal i2s_count: integer range 0 to 25;
    signal clock_12: std_logic:='0';
    signal aud_bk_counter: integer range 0 to 9:=0;
    signal reset: std_logic:='0';
    signal indexR: integer range -2 to 23:=-2; 
    signal indexL: integer range -2 to 23:=-2; 


begin 
aud_dalr<=data_clock; 
aud_data_out<=aud_out_bit;
aud_bk<=aud_bk_clock;
clock_12_out<=clock_12; 

process(master_clock)
begin
    if rising_edge(master_clock) then 
        
        -- Main Clock 12.5HZ for WM8731 (AUD_XCK)
        if(clock_12_count<1) then 
            clock_12_count <= clock_12_count +1; 
        else 
            clock_12_count<=0; 
            clock_12 <= not clock_12; 
        end if;

        -- Data Clock (DACLRC)
        if(daclrc_count<519) then 
            daclrc_count <= daclrc_count + 1; 
        else 
            daclrc_count <= 0;
            data_clock <= not data_clock;  
        end if; 

        -- Bit clock (AUD_BCLK)
        if(aud_bk_counter<9) then 
            aud_bk_counter<=aud_bk_counter+1;
        else 
            aud_bk_counter<=0;
            aud_bk_clock <= not aud_bk_clock; 
        end if; 
    end if; 
end process; 

process(data_clock, aud_bk_clock)
begin 
if (data_clock='0') then
    indexR<=-1;
elsif rising_edge(aud_bk_clock) then
    indexR <= indexR + 1;
end if;
end process;
process(data_clock, aud_bk_clock)
begin 
if (data_clock='1') then
    indexL<=-1;
elsif rising_edge(aud_bk_clock) then
    indexL <= indexL + 1;
end if;
end process;



process(data_clock, aud_bk_clock)
begin 
    if falling_edge(data_clock) then
        sample_index <= (sample_index + 1) mod ARRAY_SIZE;
    end if;
        
    if falling_edge(aud_bk_clock) then
        if (i2s_count < 1) then 
            i2s_count <= i2s_count + 1;
        elsif (i2s_count<24) then
            if (data_clock='0') then
                case keys is 
                    when "0111" =>
                        aud_out_bit <= aud_out_sample(sample_index)(indexL);
                    when "1011" => 
                        aud_out_bit <= aud_out_sample1(sample_index)(indexL);
                    when "1101" => 
                        aud_out_bit <= aud_out_sample2(sample_index)(indexL);
                    when "1110" => 
                        aud_out_bit <= aud_out_sample3(sample_index)(indexL);
                    when others =>
                        aud_out_bit<='0';
                end case;
            else
                case keys is 
                    when "0111" =>
                        aud_out_bit <= aud_out_sample(sample_index)(indexR);
                    when "1011" => 
                        aud_out_bit <= aud_out_sample1(sample_index)(indexR);
                    when "1101" => 
                        aud_out_bit <= aud_out_sample2(sample_index)(indexR);
                    when "1110" => 
                        aud_out_bit <= aud_out_sample3(sample_index)(indexR);
                    when others =>
                        aud_out_bit<='0';
                end case; 
            end if;
                i2s_count <=i2s_count + 1; 
            else
                i2s_count <=0;
        end if; 
    end if; 
end process;

end gen;
