library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity audio_gen is 
port (
    aud_clock: in std_logic;
    sw: in std_logic_vector(9 downto 0);
    ledr: OUT std_logic; 
    aud_bk: out std_logic;
    aud_dalr: out std_logic;
    aud_data: out std_logic
);
end audio_gen; 

architecture gen of audio_gen is 
    signal clk_en: std_logic:='0';
    signal send_flag: std_logic:='0';
    signal index: integer range 0 to 31:=0;
    signal sample_index: integer range 0 to 24:=0;
    signal aud_idx: std_logic := '0';
    signal aud_out: std_logic_vector(31 downto 0):=(others=>'0');
    type BinArrray is array(0 to 999) of std_logic_vector(31 downto 0);
    signal aud_out_sample: BinArrray :=( "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000"
    ,"11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000",
    "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001",
    "00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111",
    "11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111100000000","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111","11111111111111111111111111111111");
    signal aud_scale: integer range 0 to 300:=0;
    signal data_clock: std_logic:='0';
    signal aud_out_bit: std_logic;  
    constant ARRAY_SIZE: natural :=1000;
    signal bk_count: integer range 0 to 15:=0;
    signal aud_bk_clock: std_logic:='0';

begin 
aud_dalr<=data_clock; 
aud_data<=aud_out_bit;
aud_bk<=aud_bk_clock; 

process(aud_clock)
begin 
    if rising_edge(aud_clock) then
        if( aud_scale < 260) then 
            aud_scale <=aud_scale + 1; 
        else 
            data_clock <= not data_clock;
            aud_scale <=0;  
        end if;

        if (bk_count<16) then 
            bk_count<=bk_count+1;
        else
            aud_bk_clock<= not aud_bk_clock; 
            bk_count<=0;

        end if; 

    end if; 
end process;

process(data_clock)
begin 
        if rising_edge(data_clock) then
            if (index<31) then 
                aud_out_bit <= aud_out_sample(sample_index)(index);
                index <= index +1; 
            else
                aud_out_bit <= aud_out_sample(sample_index)(index);
                index <= 0;
                sample_index <= (sample_index + 1) mod ARRAY_SIZE;
            end if;
        end if; 
end process;


-- aud_bk<=aud_clock;
--     process(aud_clock)
--     begin
--         if falling_edge(aud_clock) then

--                 aud_dalr<=clk_en;
--                 if (aud_scale<250) then 
--                     aud_scale<=aud_scale+1;
--                     clk_en<='0';
--                 else 
--                     aud_scale<=0;
--                     -- aud_out<="00000000000000000111111111111111";
--                     aud_out<=aud_out_sample(sample_index);
--                     sample_index<=(sample_index+1)mod ARRAY_SIZE;
--                     clk_en<='1';
--                 end if; 

--                 if (clk_en='1') then
--                     index<=31;
--                     send_flag<='1';
--                 end if; 

--                 if (send_flag='1') then 
--                     if (index>0) then
--                         index<=index-1;
--                     else
--                         send_flag<='0';
--                     end if; 
--                     aud_data<=aud_out(index);
--                 end if;
--         end if;
--     end process;
end gen;
