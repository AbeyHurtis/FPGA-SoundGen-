library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity audio_gen is 
port (
    master_clock: in std_logic;
    clock_12_out: out std_logic:='0';
    sw: in std_logic_vector(9 downto 0);
    ledr: OUT std_logic; 
    aud_bk: out std_logic:='0';
    aud_dalr: out std_logic:='0';
    aud_data_out: out std_logic
);
end audio_gen; 

architecture gen of audio_gen is 
    signal clk_en: std_logic:='0';
    signal send_flag: std_logic:='0';
    signal index: integer range 0 to 23:=0;
    signal sample_index: integer range 0 to 23:=0;
    signal aud_idx: std_logic := '0';
    signal aud_out: std_logic_vector(23 downto 0):=(others=>'0');
    type BinArrray is array(0 to 999) of std_logic_vector(23 downto 0);
    signal aud_out_sample: BinArrray :=("000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","111111111111111100000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","111111111111111100000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111100000000",
    "000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001","000000000000000000000001",
    "000000000000000000000001","000000000000000000000001","000000000000000000000000","000000000000000000000000","000000000000000000000000","000000000000000000000000",
    "111111111111111100000000","111111111111111100000000","111111111111111100000000","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111",
    "111111111111111111111111","111111111111111111111111","111111111111111111111111","111111111111111111111111");
    signal daclrc_count: integer range 0 to 519:=0;
    signal data_clock: std_logic:='0';
    signal aud_out_bit: std_logic;  
    constant ARRAY_SIZE: natural :=1000;
    signal bk_count: integer range 0 to 15:=0;
    signal aud_bk_clock: std_logic:='0';
    signal clock_12_count: integer range 0 to 1:=0;
    signal i2s_count: integer range 0 to 25;
    signal clock_12: std_logic:='0';
    signal aud_bk_counter: integer range 0 to 9:=0;


begin 
aud_dalr<=data_clock; 
aud_data_out<=aud_out_bit;
aud_bk<=aud_bk_clock; 

process(master_clock)
begin
    if rising_edge(master_clock) then 
        
        -- Main Clock 12.5HZ for WM8731 (AUD_XCK)
        if(clock_12_count<1) then 
            clock_12_count <= clock_12_count +1; 
        else 
            clock_12_count<=0; 
            clock_12 <= not clock_12; 
        end if;

        -- Data Clock (DACLRC)
        if(daclrc_count<519) then 
            daclrc_count <= daclrc_count + 1; 
        else 
            daclrc_count <= 0;
            data_clock <= not data_clock;  
        end if; 

        -- Bit clock (AUD_BCLK)
        if(aud_bk_counter<9) then 
            aud_bk_counter<=aud_bk_counter+1;
        else 
            aud_bk_counter<=0;
            aud_bk_clock <= not aud_bk_clock; 
        end if; 
    end if; 
end process; 



process(data_clock)
begin 
    index<=0;
    if falling_edge(data_clock) then
        sample_index <= (sample_index + 1) mod ARRAY_SIZE;
    end if; 
end process;

process(aud_bk_clock)
begin 
        if falling_edge(aud_bk_clock) then 
            if (i2s_count < 1) then 
                i2s_count <= i2s_count + 1;
            elsif (i2s_count<24) then
                i2s_count <=i2s_count + 1;  
                aud_out_bit <= aud_out_sample(sample_index)(index);
            end if; 
        end if; 
end process; 
end gen;
